module main

fn main() {
    println('Hallo Welt')
}